module packed_unpacked_array;
bit  [3:0][7:0]arr[2][4];

initial begin
foreach(arr[i])begin
foreach(arr[i][j])begin
arr[i][j]=$urandom;
$display("packed & unpacked elements[%0d][%0d]:0x%0h",i,j,arr[i][j]);
$display("arr=%p",arr);
$display("arr[0][0][2]=0x%0h",arr[0][0][2]);
end
end
end
endmodule

output
 Loading work.packed_unpacked_array(fast)
run
# packed & unpacked elements[0][0]:0xce46aa23
# arr='{'{'{206, 70, 170, 35}, '{0, 0, 0, 0}, '{0, 0, 0, 0}, '{0, 0, 0, 0}}, '{'{0, 0, 0, 0}, '{0, 0, 0, 0}, '{0, 0, 0, 0}, '{0, 0, 0, 0}}}
# arr[0][0][2]=0x46
# packed & unpacked elements[0][1]:0xa01b6e32
# arr='{'{'{206, 70, 170, 35}, '{160, 27, 110, 50}, '{0, 0, 0, 0}, '{0, 0, 0, 0}}, '{'{0, 0, 0, 0}, '{0, 0, 0, 0}, '{0, 0, 0, 0}, '{0, 0, 0, 0}}}
# arr[0][0][2]=0x46
# packed & unpacked elements[0][2]:0x5cb53a0a
# arr='{'{'{206, 70, 170, 35}, '{160, 27, 110, 50}, '{92, 181, 58, 10}, '{0, 0, 0, 0}}, '{'{0, 0, 0, 0}, '{0, 0, 0, 0}, '{0, 0, 0, 0}, '{0, 0, 0, 0}}}
# arr[0][0][2]=0x46
# packed & unpacked elements[0][3]:0x8b4e9f1d
# arr='{'{'{206, 70, 170, 35}, '{160, 27, 110, 50}, '{92, 181, 58, 10}, '{139, 78, 159, 29}}, '{'{0, 0, 0, 0}, '{0, 0, 0, 0}, '{0, 0, 0, 0}, '{0, 0, 0, 0}}}
# arr[0][0][2]=0x46
# packed & unpacked elements[1][0]:0xa80385b8
# arr='{'{'{206, 70, 170, 35}, '{160, 27, 110, 50}, '{92, 181, 58, 10}, '{139, 78, 159, 29}}, '{'{168, 3, 133, 184}, '{0, 0, 0, 0}, '{0, 0, 0, 0}, '{0, 0, 0, 0}}}
# arr[0][0][2]=0x46
# packed & unpacked elements[1][1]:0x69968eda
# arr='{'{'{206, 70, 170, 35}, '{160, 27, 110, 50}, '{92, 181, 58, 10}, '{139, 78, 159, 29}}, '{'{168, 3, 133, 184}, '{105, 150, 142, 218}, '{0, 0, 0, 0}, '{0, 0, 0, 0}}}
# arr[0][0][2]=0x46
# packed & unpacked elements[1][2]:0x13c11ac0
# arr='{'{'{206, 70, 170, 35}, '{160, 27, 110, 50}, '{92, 181, 58, 10}, '{139, 78, 159, 29}}, '{'{168, 3, 133, 184}, '{105, 150, 142, 218}, '{19, 193, 26, 192}, '{0, 0, 0, 0}}}
# arr[0][0][2]=0x46
# packed & unpacked elements[1][3]:0xe0a228ac
# arr='{'{'{206, 70, 170, 35}, '{160, 27, 110, 50}, '{92, 181, 58, 10}, '{139, 78, 159, 29}}, '{'{168, 3, 133, 184}, '{105, 150, 142, 218}, '{19, 193, 26, 192}, '{224, 162, 40, 172}}}
# arr[0][0][2]=0x46
