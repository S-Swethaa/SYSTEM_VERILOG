# Loading sv_std.std
# Loading work.design_sv_unit(fast)
# Loading work.test(fast)
# Loading work.testbench(fast)
# Loading work.intf(fast__2)
# Loading work.sync_fifo(fast)
# Loading work.intf(fast)
# 
# run -all
#    Generator   
# Time=0 | w_en=0 | r_en=0 | din=bb | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=6 | w_en=0 | r_en=0 | din=0 | dataout=0 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=6 | w_en=0 | r_en=0 | din=0 | dataout=0 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=6 | w_en=0 | r_en=1 | din=e1 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=16 | w_en=0 | r_en=0 | din=0 | dataout=0 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=16 | w_en=0 | r_en=0 | din=0 | dataout=0 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=16 | w_en=1 | r_en=0 | din=81 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=25 | w_en=0 | r_en=0 | din=bb | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=26 | w_en=0 | r_en=0 | din=0 | dataout=0 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=26 | w_en=0 | r_en=0 | din=0 | dataout=0 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=26 | w_en=1 | r_en=1 | din=62 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=35 | w_en=0 | r_en=1 | din=e1 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=36 | w_en=0 | r_en=0 | din=bb | dataout=0 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=36 | w_en=0 | r_en=0 | din=bb | dataout=0 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=36 | w_en=1 | r_en=1 | din=1d | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=45 | w_en=1 | r_en=0 | din=81 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=46 | w_en=0 | r_en=0 | din=e1 | dataout=0 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=46 | w_en=0 | r_en=0 | din=e1 | dataout=0 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=46 | w_en=0 | r_en=1 | din=f7 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=55 | w_en=1 | r_en=1 | din=62 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=56 | w_en=1 | r_en=0 | din=81 | dataout=0 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=56 | w_en=1 | r_en=0 | din=81 | dataout=0 | empty=0 | full=0
# ***********************************
# Writing 81 to mem[0]
#    Generator   
# Time=56 | w_en=0 | r_en=1 | din=70 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=65 | w_en=1 | r_en=1 | din=1d | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=66 | w_en=1 | r_en=1 | din=62 | dataout=81 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=66 | w_en=1 | r_en=1 | din=62 | dataout=81 | empty=0 | full=0
# ***********************************
# Writing 62 to mem[1]
# Expecting 81 from mem[0]
# -------------------------------------------
# PASS
# -------------------------------------------
#    Generator   
# Time=66 | w_en=1 | r_en=0 | din=43 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=75 | w_en=0 | r_en=1 | din=f7 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=76 | w_en=1 | r_en=1 | din=1d | dataout=62 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=76 | w_en=1 | r_en=1 | din=1d | dataout=62 | empty=0 | full=0
# ***********************************
# Writing 1d to mem[2]
# Expecting 62 from mem[1]
# -------------------------------------------
# PASS
# -------------------------------------------
#    Generator   
# Time=76 | w_en=0 | r_en=1 | din=78 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=85 | w_en=0 | r_en=1 | din=70 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=86 | w_en=0 | r_en=1 | din=f7 | dataout=1d | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=86 | w_en=0 | r_en=1 | din=f7 | dataout=1d | empty=1 | full=0
# ***********************************
#    Generator   
# Time=86 | w_en=1 | r_en=1 | din=a1 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=95 | w_en=1 | r_en=0 | din=43 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=96 | w_en=0 | r_en=0 | din=70 | dataout=1d | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=96 | w_en=0 | r_en=0 | din=70 | dataout=1d | empty=1 | full=0
# ***********************************
#    Generator   
# Time=96 | w_en=1 | r_en=0 | din=84 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=105 | w_en=0 | r_en=1 | din=78 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=106 | w_en=1 | r_en=0 | din=43 | dataout=1d | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=106 | w_en=1 | r_en=0 | din=43 | dataout=1d | empty=0 | full=0
# ***********************************
# Writing 43 to mem[3]
#    Generator   
# Time=106 | w_en=1 | r_en=0 | din=d8 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=115 | w_en=1 | r_en=1 | din=a1 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=116 | w_en=0 | r_en=1 | din=78 | dataout=43 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=116 | w_en=0 | r_en=1 | din=78 | dataout=43 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=116 | w_en=0 | r_en=1 | din=25 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=125 | w_en=1 | r_en=0 | din=84 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=126 | w_en=1 | r_en=0 | din=a1 | dataout=43 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=126 | w_en=1 | r_en=0 | din=a1 | dataout=43 | empty=0 | full=0
# ***********************************
# Writing a1 to mem[4]
#    Generator   
# Time=126 | w_en=0 | r_en=1 | din=29 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=135 | w_en=1 | r_en=0 | din=d8 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=136 | w_en=1 | r_en=0 | din=84 | dataout=43 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=136 | w_en=1 | r_en=0 | din=84 | dataout=43 | empty=0 | full=0
# ***********************************
# Writing 84 to mem[5]
#    Generator   
# Time=136 | w_en=0 | r_en=0 | din=ab | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=145 | w_en=0 | r_en=1 | din=25 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=146 | w_en=1 | r_en=0 | din=d8 | dataout=43 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=146 | w_en=1 | r_en=0 | din=d8 | dataout=43 | empty=0 | full=0
# ***********************************
# Writing d8 to mem[6]
#    Generator   
# Time=146 | w_en=1 | r_en=1 | din=e0 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=155 | w_en=0 | r_en=1 | din=29 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=156 | w_en=0 | r_en=1 | din=25 | dataout=a1 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=156 | w_en=0 | r_en=1 | din=25 | dataout=a1 | empty=0 | full=0
# ***********************************
# Expecting 1d from mem[2]
# -------------------------------------------
# FAIL
# -------------------------------------------
#    Generator   
# Time=156 | w_en=1 | r_en=1 | din=59 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=165 | w_en=0 | r_en=0 | din=ab | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=166 | w_en=0 | r_en=1 | din=29 | dataout=84 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=166 | w_en=0 | r_en=1 | din=29 | dataout=84 | empty=0 | full=0
# ***********************************
# Expecting 43 from mem[3]
# -------------------------------------------
# FAIL
# -------------------------------------------
#    Generator   
# Time=166 | w_en=1 | r_en=1 | din=16 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=175 | w_en=1 | r_en=1 | din=e0 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=176 | w_en=0 | r_en=0 | din=ab | dataout=84 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=176 | w_en=0 | r_en=0 | din=ab | dataout=84 | empty=0 | full=0
# ***********************************
#    Generator   
# Time=176 | w_en=0 | r_en=0 | din=c1 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=185 | w_en=1 | r_en=1 | din=59 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=186 | w_en=1 | r_en=1 | din=e0 | dataout=d8 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=186 | w_en=1 | r_en=1 | din=e0 | dataout=d8 | empty=0 | full=0
# ***********************************
# Writing e0 to mem[7]
# Expecting a1 from mem[4]
# -------------------------------------------
# FAIL
# -------------------------------------------
#    Generator   
# Time=186 | w_en=0 | r_en=0 | din=5 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=195 | w_en=1 | r_en=1 | din=16 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=196 | w_en=1 | r_en=1 | din=59 | dataout=e0 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=196 | w_en=1 | r_en=1 | din=59 | dataout=e0 | empty=0 | full=0
# ***********************************
# Writing 59 to mem[8]
# Expecting 84 from mem[5]
# -------------------------------------------
# FAIL
# -------------------------------------------
#    Generator   
# Time=196 | w_en=0 | r_en=1 | din=32 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=205 | w_en=0 | r_en=0 | din=c1 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=206 | w_en=1 | r_en=1 | din=16 | dataout=59 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=206 | w_en=1 | r_en=1 | din=16 | dataout=59 | empty=0 | full=0
# ***********************************
# Writing 16 to mem[9]
# Expecting d8 from mem[6]
# -------------------------------------------
# FAIL
# -------------------------------------------
#    Generator   
# Time=206 | w_en=1 | r_en=0 | din=fb | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=215 | w_en=0 | r_en=0 | din=5 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=216 | w_en=0 | r_en=0 | din=c1 | dataout=59 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=216 | w_en=0 | r_en=0 | din=c1 | dataout=59 | empty=0 | full=0
# ***********************************
#    Generator   
# Time=216 | w_en=0 | r_en=1 | din=65 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=225 | w_en=0 | r_en=1 | din=32 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=226 | w_en=0 | r_en=0 | din=5 | dataout=59 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=226 | w_en=0 | r_en=0 | din=5 | dataout=59 | empty=0 | full=0
# ***********************************
#    Generator   
# Time=226 | w_en=1 | r_en=1 | din=a6 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=235 | w_en=1 | r_en=0 | din=fb | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=236 | w_en=0 | r_en=1 | din=32 | dataout=16 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=236 | w_en=0 | r_en=1 | din=32 | dataout=16 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=236 | w_en=0 | r_en=1 | din=49 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=245 | w_en=0 | r_en=1 | din=65 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=246 | w_en=1 | r_en=0 | din=fb | dataout=16 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=246 | w_en=1 | r_en=0 | din=fb | dataout=16 | empty=0 | full=0
# ***********************************
# Writing fb to mem[10]
#    Generator   
# Time=246 | w_en=0 | r_en=1 | din=e6 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=255 | w_en=1 | r_en=1 | din=a6 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=256 | w_en=0 | r_en=1 | din=65 | dataout=fb | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=256 | w_en=0 | r_en=1 | din=65 | dataout=fb | empty=1 | full=0
# ***********************************
#    Generator   
# Time=256 | w_en=1 | r_en=1 | din=d7 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=265 | w_en=0 | r_en=1 | din=49 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=266 | w_en=1 | r_en=0 | din=a6 | dataout=fb | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=266 | w_en=1 | r_en=0 | din=a6 | dataout=fb | empty=0 | full=0
# ***********************************
# Writing a6 to mem[11]
#    Generator   
# Time=266 | w_en=1 | r_en=1 | din=2d | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=275 | w_en=0 | r_en=1 | din=e6 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=276 | w_en=0 | r_en=1 | din=49 | dataout=a6 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=276 | w_en=0 | r_en=1 | din=49 | dataout=a6 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=276 | w_en=0 | r_en=1 | din=bf | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=285 | w_en=1 | r_en=1 | din=d7 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=286 | w_en=0 | r_en=0 | din=e6 | dataout=a6 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=286 | w_en=0 | r_en=0 | din=e6 | dataout=a6 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=286 | w_en=0 | r_en=1 | din=38 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=295 | w_en=1 | r_en=1 | din=2d | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=296 | w_en=1 | r_en=0 | din=d7 | dataout=a6 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=296 | w_en=1 | r_en=0 | din=d7 | dataout=a6 | empty=0 | full=0
# ***********************************
# Writing d7 to mem[12]
#    Generator   
# Time=296 | w_en=1 | r_en=0 | din=6a | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=305 | w_en=0 | r_en=1 | din=bf | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=306 | w_en=1 | r_en=1 | din=2d | dataout=d7 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=306 | w_en=1 | r_en=1 | din=2d | dataout=d7 | empty=0 | full=0
# ***********************************
# Writing 2d to mem[13]
# Expecting e0 from mem[7]
# -------------------------------------------
# FAIL
# -------------------------------------------
#    Generator   
# Time=306 | w_en=0 | r_en=0 | din=94 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=315 | w_en=0 | r_en=1 | din=38 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=316 | w_en=0 | r_en=1 | din=bf | dataout=2d | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=316 | w_en=0 | r_en=1 | din=bf | dataout=2d | empty=1 | full=0
# ***********************************
#    Generator   
# Time=316 | w_en=0 | r_en=1 | din=d1 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=325 | w_en=1 | r_en=0 | din=6a | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=326 | w_en=0 | r_en=0 | din=38 | dataout=2d | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=326 | w_en=0 | r_en=0 | din=38 | dataout=2d | empty=1 | full=0
# ***********************************
#    Generator   
# Time=326 | w_en=0 | r_en=0 | din=7b | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=335 | w_en=0 | r_en=0 | din=94 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=336 | w_en=1 | r_en=0 | din=6a | dataout=2d | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=336 | w_en=1 | r_en=0 | din=6a | dataout=2d | empty=0 | full=0
# ***********************************
# Writing 6a to mem[14]
#    Generator   
# Time=336 | w_en=1 | r_en=1 | din=ad | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=345 | w_en=0 | r_en=1 | din=d1 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=346 | w_en=0 | r_en=0 | din=94 | dataout=2d | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=346 | w_en=0 | r_en=0 | din=94 | dataout=2d | empty=0 | full=0
# ***********************************
#    Generator   
# Time=346 | w_en=0 | r_en=0 | din=85 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=355 | w_en=0 | r_en=0 | din=7b | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=356 | w_en=0 | r_en=1 | din=d1 | dataout=6a | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=356 | w_en=0 | r_en=1 | din=d1 | dataout=6a | empty=1 | full=0
# ***********************************
#    Generator   
# Time=356 | w_en=1 | r_en=1 | din=8 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=365 | w_en=1 | r_en=1 | din=ad | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=366 | w_en=0 | r_en=0 | din=7b | dataout=6a | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=366 | w_en=0 | r_en=0 | din=7b | dataout=6a | empty=1 | full=0
# ***********************************
#    Generator   
# Time=366 | w_en=0 | r_en=1 | din=56 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=375 | w_en=0 | r_en=0 | din=85 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=376 | w_en=1 | r_en=0 | din=ad | dataout=6a | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=376 | w_en=1 | r_en=0 | din=ad | dataout=6a | empty=0 | full=0
# ***********************************
# Writing ad to mem[15]
#    Generator   
# Time=376 | w_en=1 | r_en=0 | din=dc | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=385 | w_en=1 | r_en=1 | din=8 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=386 | w_en=0 | r_en=0 | din=85 | dataout=6a | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=386 | w_en=0 | r_en=0 | din=85 | dataout=6a | empty=0 | full=0
# ***********************************
#    Generator   
# Time=386 | w_en=0 | r_en=1 | din=76 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=395 | w_en=0 | r_en=1 | din=56 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=396 | w_en=1 | r_en=1 | din=8 | dataout=ad | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=396 | w_en=1 | r_en=1 | din=8 | dataout=ad | empty=0 | full=0
# ***********************************
# Writing 8 to mem[0]
# Expecting 59 from mem[8]
# -------------------------------------------
# FAIL
# -------------------------------------------
#    Generator   
# Time=396 | w_en=1 | r_en=0 | din=72 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=405 | w_en=1 | r_en=0 | din=dc | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=406 | w_en=0 | r_en=1 | din=56 | dataout=8 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=406 | w_en=0 | r_en=1 | din=56 | dataout=8 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=406 | w_en=0 | r_en=0 | din=97 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=415 | w_en=0 | r_en=1 | din=76 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=416 | w_en=1 | r_en=0 | din=dc | dataout=8 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=416 | w_en=1 | r_en=0 | din=dc | dataout=8 | empty=0 | full=0
# ***********************************
# Writing dc to mem[1]
#    Generator   
# Time=416 | w_en=1 | r_en=0 | din=e | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=425 | w_en=1 | r_en=0 | din=72 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=426 | w_en=0 | r_en=1 | din=76 | dataout=dc | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=426 | w_en=0 | r_en=1 | din=76 | dataout=dc | empty=1 | full=0
# ***********************************
#    Generator   
# Time=426 | w_en=0 | r_en=0 | din=b2 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=435 | w_en=0 | r_en=0 | din=97 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=436 | w_en=1 | r_en=0 | din=72 | dataout=dc | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=436 | w_en=1 | r_en=0 | din=72 | dataout=dc | empty=0 | full=0
# ***********************************
# Writing 72 to mem[2]
#    Generator   
# Time=436 | w_en=1 | r_en=1 | din=48 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=445 | w_en=1 | r_en=0 | din=e | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=446 | w_en=0 | r_en=0 | din=97 | dataout=dc | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=446 | w_en=0 | r_en=0 | din=97 | dataout=dc | empty=0 | full=0
# ***********************************
#    Generator   
# Time=446 | w_en=0 | r_en=1 | din=e | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=455 | w_en=0 | r_en=0 | din=b2 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=456 | w_en=1 | r_en=0 | din=e | dataout=dc | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=456 | w_en=1 | r_en=0 | din=e | dataout=dc | empty=0 | full=0
# ***********************************
# Writing e to mem[3]
#    Generator   
# Time=456 | w_en=0 | r_en=0 | din=65 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=465 | w_en=1 | r_en=1 | din=48 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=466 | w_en=0 | r_en=0 | din=b2 | dataout=dc | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=466 | w_en=0 | r_en=0 | din=b2 | dataout=dc | empty=0 | full=0
# ***********************************
#    Generator   
# Time=466 | w_en=0 | r_en=1 | din=43 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=475 | w_en=0 | r_en=1 | din=e | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=476 | w_en=1 | r_en=1 | din=48 | dataout=72 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=476 | w_en=1 | r_en=1 | din=48 | dataout=72 | empty=0 | full=0
# ***********************************
# Writing 48 to mem[4]
# Expecting 16 from mem[9]
# -------------------------------------------
# FAIL
# -------------------------------------------
#    Generator   
# Time=476 | w_en=0 | r_en=1 | din=76 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=485 | w_en=0 | r_en=0 | din=65 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=486 | w_en=0 | r_en=1 | din=e | dataout=e | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=486 | w_en=0 | r_en=1 | din=e | dataout=e | empty=0 | full=0
# ***********************************
# Expecting fb from mem[10]
# -------------------------------------------
# FAIL
# -------------------------------------------
#    Generator   
# Time=486 | w_en=0 | r_en=0 | din=95 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=495 | w_en=0 | r_en=1 | din=43 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=496 | w_en=0 | r_en=0 | din=65 | dataout=e | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=496 | w_en=0 | r_en=0 | din=65 | dataout=e | empty=0 | full=0
# ***********************************
#    Generator   
# Time=496 | w_en=1 | r_en=1 | din=40 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=505 | w_en=0 | r_en=1 | din=76 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=506 | w_en=0 | r_en=1 | din=43 | dataout=48 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=506 | w_en=0 | r_en=1 | din=43 | dataout=48 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=506 | w_en=1 | r_en=1 | din=a5 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=515 | w_en=0 | r_en=0 | din=95 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=516 | w_en=0 | r_en=0 | din=76 | dataout=48 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=516 | w_en=0 | r_en=0 | din=76 | dataout=48 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=516 | w_en=1 | r_en=1 | din=96 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=525 | w_en=1 | r_en=1 | din=40 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=526 | w_en=0 | r_en=0 | din=95 | dataout=48 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=526 | w_en=0 | r_en=0 | din=95 | dataout=48 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=526 | w_en=1 | r_en=0 | din=93 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=535 | w_en=1 | r_en=1 | din=a5 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=536 | w_en=1 | r_en=0 | din=40 | dataout=48 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=536 | w_en=1 | r_en=0 | din=40 | dataout=48 | empty=0 | full=0
# ***********************************
# Writing 40 to mem[5]
#    Generator   
# Time=536 | w_en=0 | r_en=1 | din=69 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=545 | w_en=1 | r_en=1 | din=96 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=546 | w_en=1 | r_en=1 | din=a5 | dataout=40 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=546 | w_en=1 | r_en=1 | din=a5 | dataout=40 | empty=0 | full=0
# ***********************************
# Writing a5 to mem[6]
# Expecting a6 from mem[11]
# -------------------------------------------
# FAIL
# -------------------------------------------
#    Generator   
# Time=546 | w_en=0 | r_en=1 | din=42 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=555 | w_en=1 | r_en=0 | din=93 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=556 | w_en=1 | r_en=1 | din=96 | dataout=a5 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=556 | w_en=1 | r_en=1 | din=96 | dataout=a5 | empty=0 | full=0
# ***********************************
# Writing 96 to mem[7]
# Expecting d7 from mem[12]
# -------------------------------------------
# FAIL
# -------------------------------------------
#    Generator   
# Time=556 | w_en=0 | r_en=1 | din=4e | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=565 | w_en=0 | r_en=1 | din=69 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=566 | w_en=1 | r_en=0 | din=93 | dataout=a5 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=566 | w_en=1 | r_en=0 | din=93 | dataout=a5 | empty=0 | full=0
# ***********************************
# Writing 93 to mem[8]
#    Generator   
# Time=566 | w_en=1 | r_en=0 | din=6c | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=575 | w_en=0 | r_en=1 | din=42 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=576 | w_en=0 | r_en=1 | din=69 | dataout=96 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=576 | w_en=0 | r_en=1 | din=69 | dataout=96 | empty=0 | full=0
# ***********************************
# Expecting 2d from mem[13]
# -------------------------------------------
# FAIL
# -------------------------------------------
#    Generator   
# Time=576 | w_en=1 | r_en=1 | din=92 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=585 | w_en=0 | r_en=1 | din=4e | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=586 | w_en=0 | r_en=1 | din=42 | dataout=93 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=586 | w_en=0 | r_en=1 | din=42 | dataout=93 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=586 | w_en=0 | r_en=1 | din=2f | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=595 | w_en=1 | r_en=0 | din=6c | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=596 | w_en=0 | r_en=0 | din=4e | dataout=93 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=596 | w_en=0 | r_en=0 | din=4e | dataout=93 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=596 | w_en=1 | r_en=0 | din=9c | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=605 | w_en=1 | r_en=1 | din=92 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=606 | w_en=1 | r_en=0 | din=6c | dataout=93 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=606 | w_en=1 | r_en=0 | din=6c | dataout=93 | empty=0 | full=0
# ***********************************
# Writing 6c to mem[9]
#    Generator   
# Time=606 | w_en=0 | r_en=1 | din=95 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=615 | w_en=0 | r_en=1 | din=2f | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=616 | w_en=1 | r_en=1 | din=92 | dataout=6c | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=616 | w_en=1 | r_en=1 | din=92 | dataout=6c | empty=0 | full=0
# ***********************************
# Writing 92 to mem[10]
# Expecting 6a from mem[14]
# -------------------------------------------
# FAIL
# -------------------------------------------
#    Generator   
# Time=616 | w_en=0 | r_en=1 | din=1 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=625 | w_en=1 | r_en=0 | din=9c | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=626 | w_en=0 | r_en=1 | din=2f | dataout=92 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=626 | w_en=0 | r_en=1 | din=2f | dataout=92 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=626 | w_en=0 | r_en=1 | din=56 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=635 | w_en=0 | r_en=1 | din=95 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=636 | w_en=1 | r_en=0 | din=9c | dataout=92 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=636 | w_en=1 | r_en=0 | din=9c | dataout=92 | empty=0 | full=0
# ***********************************
# Writing 9c to mem[11]
#    Generator   
# Time=636 | w_en=1 | r_en=0 | din=eb | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=645 | w_en=0 | r_en=1 | din=1 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=646 | w_en=0 | r_en=1 | din=95 | dataout=9c | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=646 | w_en=0 | r_en=1 | din=95 | dataout=9c | empty=1 | full=0
# ***********************************
#    Generator   
# Time=646 | w_en=0 | r_en=0 | din=1c | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=655 | w_en=0 | r_en=1 | din=56 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=656 | w_en=0 | r_en=0 | din=1 | dataout=9c | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=656 | w_en=0 | r_en=0 | din=1 | dataout=9c | empty=1 | full=0
# ***********************************
#    Generator   
# Time=656 | w_en=1 | r_en=1 | din=78 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=665 | w_en=1 | r_en=0 | din=eb | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=666 | w_en=0 | r_en=0 | din=56 | dataout=9c | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=666 | w_en=0 | r_en=0 | din=56 | dataout=9c | empty=1 | full=0
# ***********************************
#    Generator   
# Time=666 | w_en=0 | r_en=1 | din=cf | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=675 | w_en=0 | r_en=0 | din=1c | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=676 | w_en=1 | r_en=0 | din=eb | dataout=9c | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=676 | w_en=1 | r_en=0 | din=eb | dataout=9c | empty=0 | full=0
# ***********************************
# Writing eb to mem[12]
#    Generator   
# Time=676 | w_en=1 | r_en=1 | din=c7 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=685 | w_en=1 | r_en=1 | din=78 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=686 | w_en=0 | r_en=0 | din=1c | dataout=9c | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=686 | w_en=0 | r_en=0 | din=1c | dataout=9c | empty=0 | full=0
# ***********************************
#    Generator   
# Time=686 | w_en=0 | r_en=1 | din=7b | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=695 | w_en=0 | r_en=1 | din=cf | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=696 | w_en=1 | r_en=1 | din=78 | dataout=eb | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=696 | w_en=1 | r_en=1 | din=78 | dataout=eb | empty=0 | full=0
# ***********************************
# Writing 78 to mem[13]
# Expecting ad from mem[15]
# -------------------------------------------
# FAIL
# -------------------------------------------
#    Generator   
# Time=696 | w_en=0 | r_en=1 | din=5c | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=705 | w_en=1 | r_en=1 | din=c7 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=706 | w_en=0 | r_en=1 | din=cf | dataout=78 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=706 | w_en=0 | r_en=1 | din=cf | dataout=78 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=706 | w_en=1 | r_en=1 | din=28 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=715 | w_en=0 | r_en=1 | din=7b | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=716 | w_en=1 | r_en=0 | din=c7 | dataout=78 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=716 | w_en=1 | r_en=0 | din=c7 | dataout=78 | empty=0 | full=0
# ***********************************
# Writing c7 to mem[14]
#    Generator   
# Time=716 | w_en=1 | r_en=0 | din=81 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=725 | w_en=0 | r_en=1 | din=5c | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=726 | w_en=0 | r_en=1 | din=7b | dataout=c7 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=726 | w_en=0 | r_en=1 | din=7b | dataout=c7 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=726 | w_en=1 | r_en=1 | din=dd | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=735 | w_en=1 | r_en=1 | din=28 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=736 | w_en=0 | r_en=0 | din=5c | dataout=c7 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=736 | w_en=0 | r_en=0 | din=5c | dataout=c7 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=736 | w_en=0 | r_en=1 | din=b1 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=745 | w_en=1 | r_en=0 | din=81 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=746 | w_en=1 | r_en=0 | din=28 | dataout=c7 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=746 | w_en=1 | r_en=0 | din=28 | dataout=c7 | empty=0 | full=0
# ***********************************
# Writing 28 to mem[15]
#    Generator   
# Time=746 | w_en=1 | r_en=0 | din=ae | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=755 | w_en=1 | r_en=1 | din=dd | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=756 | w_en=1 | r_en=0 | din=81 | dataout=c7 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=756 | w_en=1 | r_en=0 | din=81 | dataout=c7 | empty=0 | full=0
# ***********************************
# Writing 81 to mem[0]
#    Generator   
# Time=756 | w_en=0 | r_en=1 | din=c2 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=765 | w_en=0 | r_en=1 | din=b1 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=766 | w_en=1 | r_en=1 | din=dd | dataout=28 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=766 | w_en=1 | r_en=1 | din=dd | dataout=28 | empty=0 | full=0
# ***********************************
# Writing dd to mem[1]
# Expecting 81 from mem[0]
# -------------------------------------------
# FAIL
# -------------------------------------------
#    Generator   
# Time=766 | w_en=1 | r_en=0 | din=38 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=775 | w_en=1 | r_en=0 | din=ae | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=776 | w_en=0 | r_en=1 | din=b1 | dataout=81 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=776 | w_en=0 | r_en=1 | din=b1 | dataout=81 | empty=0 | full=0
# ***********************************
# Expecting dd from mem[1]
# -------------------------------------------
# FAIL
# -------------------------------------------
#    Generator   
# Time=776 | w_en=0 | r_en=0 | din=c8 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=785 | w_en=0 | r_en=1 | din=c2 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=786 | w_en=1 | r_en=0 | din=ae | dataout=81 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=786 | w_en=1 | r_en=0 | din=ae | dataout=81 | empty=0 | full=0
# ***********************************
# Writing ae to mem[2]
#    Generator   
# Time=786 | w_en=0 | r_en=0 | din=87 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=795 | w_en=1 | r_en=0 | din=38 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=796 | w_en=0 | r_en=1 | din=c2 | dataout=dd | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=796 | w_en=0 | r_en=1 | din=c2 | dataout=dd | empty=0 | full=0
# ***********************************
# Expecting ae from mem[2]
# -------------------------------------------
# FAIL
# -------------------------------------------
#    Generator   
# Time=796 | w_en=0 | r_en=1 | din=c0 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=805 | w_en=0 | r_en=0 | din=c8 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=806 | w_en=1 | r_en=0 | din=38 | dataout=dd | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=806 | w_en=1 | r_en=0 | din=38 | dataout=dd | empty=0 | full=0
# ***********************************
# Writing 38 to mem[3]
#    Generator   
# Time=806 | w_en=0 | r_en=1 | din=b9 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=815 | w_en=0 | r_en=0 | din=87 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=816 | w_en=0 | r_en=0 | din=c8 | dataout=dd | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=816 | w_en=0 | r_en=0 | din=c8 | dataout=dd | empty=0 | full=0
# ***********************************
#    Generator   
# Time=816 | w_en=0 | r_en=0 | din=5b | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=825 | w_en=0 | r_en=1 | din=c0 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=826 | w_en=0 | r_en=0 | din=87 | dataout=dd | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=826 | w_en=0 | r_en=0 | din=87 | dataout=dd | empty=0 | full=0
# ***********************************
#    Generator   
# Time=826 | w_en=0 | r_en=0 | din=e9 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=835 | w_en=0 | r_en=1 | din=b9 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=836 | w_en=0 | r_en=1 | din=c0 | dataout=ae | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=836 | w_en=0 | r_en=1 | din=c0 | dataout=ae | empty=0 | full=0
# ***********************************
# Expecting 38 from mem[3]
# -------------------------------------------
# FAIL
# -------------------------------------------
#    Generator   
# Time=836 | w_en=1 | r_en=1 | din=52 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=845 | w_en=0 | r_en=0 | din=5b | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=846 | w_en=0 | r_en=1 | din=b9 | dataout=38 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=846 | w_en=0 | r_en=1 | din=b9 | dataout=38 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=846 | w_en=1 | r_en=1 | din=46 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=855 | w_en=0 | r_en=0 | din=e9 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=856 | w_en=0 | r_en=0 | din=5b | dataout=38 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=856 | w_en=0 | r_en=0 | din=5b | dataout=38 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=856 | w_en=0 | r_en=1 | din=a6 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=865 | w_en=1 | r_en=1 | din=52 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=866 | w_en=0 | r_en=0 | din=e9 | dataout=38 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=866 | w_en=0 | r_en=0 | din=e9 | dataout=38 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=866 | w_en=1 | r_en=1 | din=8c | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=875 | w_en=1 | r_en=1 | din=46 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=876 | w_en=1 | r_en=0 | din=52 | dataout=38 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=876 | w_en=1 | r_en=0 | din=52 | dataout=38 | empty=0 | full=0
# ***********************************
# Writing 52 to mem[4]
#    Generator   
# Time=876 | w_en=0 | r_en=1 | din=6a | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=885 | w_en=0 | r_en=1 | din=a6 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=886 | w_en=1 | r_en=1 | din=46 | dataout=52 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=886 | w_en=1 | r_en=1 | din=46 | dataout=52 | empty=0 | full=0
# ***********************************
# Writing 46 to mem[5]
# Expecting 52 from mem[4]
# -------------------------------------------
# PASS
# -------------------------------------------
#    Generator   
# Time=886 | w_en=1 | r_en=0 | din=20 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=895 | w_en=1 | r_en=1 | din=8c | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=896 | w_en=0 | r_en=1 | din=a6 | dataout=46 | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=896 | w_en=0 | r_en=1 | din=a6 | dataout=46 | empty=1 | full=0
# ***********************************
#    Generator   
# Time=896 | w_en=1 | r_en=0 | din=32 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=905 | w_en=0 | r_en=1 | din=6a | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=906 | w_en=1 | r_en=0 | din=8c | dataout=46 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=906 | w_en=1 | r_en=0 | din=8c | dataout=46 | empty=0 | full=0
# ***********************************
# Writing 8c to mem[6]
#    Generator   
# Time=906 | w_en=1 | r_en=0 | din=95 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=915 | w_en=1 | r_en=0 | din=20 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=916 | w_en=0 | r_en=1 | din=6a | dataout=8c | empty=1 | full=0
# ***********************************
#    Scoreboard   
# Time=916 | w_en=0 | r_en=1 | din=6a | dataout=8c | empty=1 | full=0
# ***********************************
#    Generator   
# Time=916 | w_en=1 | r_en=0 | din=f4 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=925 | w_en=1 | r_en=0 | din=32 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=926 | w_en=1 | r_en=0 | din=20 | dataout=8c | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=926 | w_en=1 | r_en=0 | din=20 | dataout=8c | empty=0 | full=0
# ***********************************
# Writing 20 to mem[7]
#    Generator   
# Time=926 | w_en=1 | r_en=0 | din=86 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=935 | w_en=1 | r_en=0 | din=95 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=936 | w_en=1 | r_en=0 | din=32 | dataout=8c | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=936 | w_en=1 | r_en=0 | din=32 | dataout=8c | empty=0 | full=0
# ***********************************
# Writing 32 to mem[8]
#    Generator   
# Time=936 | w_en=1 | r_en=0 | din=71 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=945 | w_en=1 | r_en=0 | din=f4 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=946 | w_en=1 | r_en=0 | din=95 | dataout=8c | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=946 | w_en=1 | r_en=0 | din=95 | dataout=8c | empty=0 | full=0
# ***********************************
# Writing 95 to mem[9]
#    Generator   
# Time=946 | w_en=0 | r_en=0 | din=63 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=955 | w_en=1 | r_en=0 | din=86 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=956 | w_en=1 | r_en=0 | din=f4 | dataout=8c | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=956 | w_en=1 | r_en=0 | din=f4 | dataout=8c | empty=0 | full=0
# ***********************************
# Writing f4 to mem[10]
#    Generator   
# Time=956 | w_en=1 | r_en=1 | din=dc | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=965 | w_en=1 | r_en=0 | din=71 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=966 | w_en=1 | r_en=0 | din=86 | dataout=8c | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=966 | w_en=1 | r_en=0 | din=86 | dataout=8c | empty=0 | full=0
# ***********************************
# Writing 86 to mem[11]
#    Generator   
# Time=966 | w_en=0 | r_en=0 | din=f2 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=975 | w_en=0 | r_en=0 | din=63 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=976 | w_en=1 | r_en=0 | din=71 | dataout=8c | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=976 | w_en=1 | r_en=0 | din=71 | dataout=8c | empty=0 | full=0
# ***********************************
# Writing 71 to mem[12]
#    Generator   
# Time=976 | w_en=0 | r_en=0 | din=63 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=985 | w_en=1 | r_en=1 | din=dc | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=986 | w_en=0 | r_en=0 | din=63 | dataout=8c | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=986 | w_en=0 | r_en=0 | din=63 | dataout=8c | empty=0 | full=0
# ***********************************
#    Generator   
# Time=986 | w_en=0 | r_en=1 | din=a6 | dataout=0 | empty=0 | full=0
# ***********************************
#    Driver   
# Time=995 | w_en=0 | r_en=0 | din=f2 | dataout=0 | empty=0 | full=0
# ***********************************
#    Monitor   
# Time=996 | w_en=1 | r_en=1 | din=dc | dataout=20 | empty=0 | full=0
# ***********************************
#    Scoreboard   
# Time=996 | w_en=1 | r_en=1 | din=dc | dataout=20 | empty=0 | full=0
# ***********************************
# Writing dc to mem[13]
# Expecting 46 from mem[5]
# -------------------------------------------
# FAIL
# -------------------------------------------
#    Generator   
# Time=996 | w_en=0 | r_en=0 | din=91 | dataout=0 | empty=0 | full=0
# ***********************************
# ** Note: $finish    : testbench.sv(41)
#    Time: 1 us  Iteration: 0  Instance: /testbench
# End time: 10:38:59 on Nov 02,2025, Elapsed time: 0:00:01
# Errors: 0, Warnings: 0
End time: 10:38:59 on Nov 02,2025, Elapsed time: 0:00:02
*** Summary *********************************************
    qrun: Errors:   0, Warnings:   0
    vlog: Errors:   0, Warnings:   0
    vopt: Errors:   0, Warnings:   1
    vsim: Errors:   0, Warnings:   0
  Totals: Errors:   0, Warnings:   1
