# Loading sv_std.std
# Loading work.design_sv_unit(fast)
# Loading work.testbench(fast)
# Loading work.intf(fast__2)
# Loading work.test(fast)
# Loading work.d_ff(fast)
# Loading work.intf(fast)
# 
# run -all
# ---- generator class signals ----
# $time=0,d=1,rst=1,q=0
# .........*..........
# ---- generator class signals ----
# $time=0,d=0,rst=0,q=0
# .........*..........
# ---- generator class signals ----
# $time=0,d=1,rst=0,q=0
# .........*..........
# ---- generator class signals ----
# $time=0,d=0,rst=1,q=0
# .........*..........
# ---- generator class signals ----
# $time=0,d=0,rst=0,q=0
# .........*..........
# ---- generator class signals ----
# $time=0,d=0,rst=0,q=0
# .........*..........
# ---- generator class signals ----
# $time=0,d=1,rst=1,q=0
# .........*..........
# ---- generator class signals ----
# $time=0,d=0,rst=0,q=0
# .........*..........
# ---- generator class signals ----
# $time=0,d=0,rst=0,q=0
# .........*..........
# ---- generator class signals ----
# $time=0,d=0,rst=1,q=0
# .........*..........
# monitor class signals
# ---- scoreboard class signal ----
# $time=6,d=0,rst=0,q=0
# .........*..........
# ***PASS***Exp=0, dut_out=0
# .....transaction done.....
# ====================================
# ---- driver class signal ----
# $time=15,d=1,rst=1,q=0
# .........*..........
# monitor class signals
# ---- scoreboard class signal ----
# $time=16,d=1,rst=1,q=0
# .........*..........
# ***PASS***Exp=0, dut_out=0
# .....transaction done.....
# ====================================
# ---- driver class signal ----
# $time=25,d=0,rst=0,q=0
# .........*..........
# monitor class signals
# ---- scoreboard class signal ----
# $time=26,d=0,rst=0,q=0
# .........*..........
# ***PASS***Exp=0, dut_out=0
# .....transaction done.....
# ====================================
# ---- driver class signal ----
# $time=35,d=1,rst=0,q=0
# .........*..........
# monitor class signals
# ---- scoreboard class signal ----
# $time=36,d=1,rst=0,q=1
# .........*..........
# ***PASS***Exp=1, dut_out=1
# .....transaction done.....
# ====================================
# ---- driver class signal ----
# $time=45,d=0,rst=1,q=0
# .........*..........
# monitor class signals
# ---- scoreboard class signal ----
# $time=46,d=0,rst=1,q=0
# .........*..........
# ***PASS***Exp=0, dut_out=0
# .....transaction done.....
# ====================================
# ---- driver class signal ----
# $time=55,d=0,rst=0,q=0
# .........*..........
# monitor class signals
# ---- scoreboard class signal ----
# $time=56,d=0,rst=0,q=0
# .........*..........
# ***PASS***Exp=0, dut_out=0
# .....transaction done.....
# ====================================
# ---- driver class signal ----
# $time=65,d=0,rst=0,q=0
# .........*..........
# monitor class signals
# ---- scoreboard class signal ----
# $time=66,d=0,rst=0,q=0
# .........*..........
# ***PASS***Exp=0, dut_out=0
# .....transaction done.....
# ====================================
# ---- driver class signal ----
# $time=75,d=1,rst=1,q=0
# .........*..........
# monitor class signals
# ---- scoreboard class signal ----
# $time=76,d=1,rst=1,q=0
# .........*..........
# ***PASS***Exp=0, dut_out=0
# .....transaction done.....
# ====================================
# ---- driver class signal ----
# $time=85,d=0,rst=0,q=0
# .........*..........
# monitor class signals
# ---- scoreboard class signal ----
# $time=86,d=0,rst=0,q=0
# .........*..........
# ***PASS***Exp=0, dut_out=0
# .....transaction done.....
# ====================================
# ---- driver class signal ----
# $time=95,d=0,rst=0,q=0
# .........*..........
# monitor class signals
# ---- scoreboard class signal ----
# $time=96,d=0,rst=0,q=0
# .........*..........
# ***PASS***Exp=0, dut_out=0
# .....transaction done.....
# ====================================
# ---- driver class signal ----
# $time=105,d=0,rst=1,q=0
# .........*..........
# ** Note: implicit $finish from program    : transaction.sv(9)
#    Time: 105 ns  Iteration: 1  Instance: /testbench/t
# End time: 09:21:44 on Oct 30,2025, Elapsed time: 0:00:01
# Errors: 0, Warnings: 0
End time: 09:21:44 on Oct 30,2025, Elapsed time: 0:00:02
*** Summary *********************************************
    qrun: Errors:   0, Warnings:   0
    vlog: Errors:   0, Warnings:   1
    vopt: Errors:   0, Warnings:   2
    vsim: Errors:   0, Warnings:   0
  Totals: Errors:   0, Warnings:   3
Finding VCD file...
./dump.vcd
