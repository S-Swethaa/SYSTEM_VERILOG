//INTERFACE
interface intf();
  logic a, b, c;
  logic sum, carry;
endinterface
