module unique_02();
 //An error warning Example
//None of if conditions are true or there is no ?else? statement
  int a;
  int b;
  
  initial begin
  a=20;
  b=30;
  unique if (a>b)
  $display("a is greater than b");
  else if (b >50)
  $display("b is greater than 50");
  else
  $display("a is equal to b");
  end

endmodule

output
Warning: unique condition not matched — no branch taken



