module packed_array_static;
bit [7:0]arr;

initial begin
arr=$urandom;
//foreach (arr[i])begin
$display("static packed_array=%b",arr);
//end
end
endmodule

output
# static packed_array=00100011
