module else_if_stmt;
int a,b;

initial begin
a=$urandom;
b=25;

if(a>b)
$display("a is greater than b",a,b);
else if(a<b)
$display("a is less than b",a,b);
else 
$display("a is equal to b",a,b);
end
endmodule

output
# a is less than b -834229725         25
